-- Copyright (C) 1991-2012 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 12.1 Build 177 11/07/2012 SJ Web Edition
-- Created on Sat May 18 16:58:07 2019

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Crazy_Machine IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
		  Ppad1_I : IN STD_LOGIC := '0';
        Ppad2_I : IN STD_LOGIC := '0';
        Ppad3_I : IN STD_LOGIC := '0';
		  Button_1 : IN STD_LOGIC := '0';
        sw9 : IN STD_LOGIC := '0';
        sw8 : IN STD_LOGIC := '0';
        led9 : OUT STD_LOGIC;
        led8 : OUT STD_LOGIC;
        led7 : OUT STD_LOGIC;
        led6 : OUT STD_LOGIC;
        led5 : OUT STD_LOGIC;
        led4 : OUT STD_LOGIC;
        StateBit_1 : OUT STD_LOGIC;
        StateBit_2 : OUT STD_LOGIC;
        StateBit_3 : OUT STD_LOGIC;
        servo1: OUT STD_LOGIC;
		  servo2: OUT STD_LOGIC;
		  servo3: OUT STD_LOGIC;
		  servo4: OUT STD_LOGIC
    );
END Crazy_Machine;

ARCHITECTURE BEHAVIOR OF Crazy_Machine IS
	 COMPONENT Timer
		PORT(
			clk     : in std_logic;
			reset    : in std_logic; -- Negative reset
			Millis : inout integer;
			Seconds : inout integer;
			Minutes : inout integer
		);
end COMPONENT;

	 COMPONENT TimerAlt
		PORT(
			clk     : in std_logic;
			reset    : in std_logic; -- Negative reset
			Millis : inout integer;
			Seconds : inout integer;
			Minutes : inout integer
		);
end COMPONENT;
    
    COMPONENT servo_pwm1
        PORT (
            clk   : IN  STD_LOGIC;
            reset : IN  STD_LOGIC;
            pos1   : IN INTEGER range 0 to 360;
            servo1 : OUT STD_LOGIC
        );
    END COMPONENT;
	 
	 COMPONENT servo_pwm2
        PORT (
            clk   : IN  STD_LOGIC;
            reset : IN  STD_LOGIC;
            pos2   : IN INTEGER range 0 to 360;
            servo2 : OUT STD_LOGIC
        );
    END COMPONENT;
	 
	 COMPONENT servo_pwm3
        PORT (
            clk   : IN  STD_LOGIC;
            reset : IN  STD_LOGIC;
            pos3   : IN INTEGER range 0 to 360;
            servo3 : OUT STD_LOGIC
        );
    END COMPONENT;
	 
	 COMPONENT servo_pwm4
        PORT (
            clk   : IN  STD_LOGIC;
            reset : IN  STD_LOGIC;
            pos4   : IN INTEGER range 0 to 360;
            servo4 : OUT STD_LOGIC
        );
    END COMPONENT;
	 
	 signal clk_out : STD_LOGIC := '0';
    TYPE type_fstate IS (State000,State001,State010,State011,State100,State101);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
	 SIGNAL pos1 : INTEGER range 0 to 360;
	 SIGNAL pos2 : INTEGER range 0 to 360;
	 SIGNAL pos3 : INTEGER range 0 to 360;
	 SIGNAL pos4 : INTEGER range 0 to 360;
	 SIGNAL Millis : INTEGER;
	 SIGNAL Seconds : INTEGER;
	 SIGNAL Minutes : INTEGER;
	 SIGNAL started : STD_LOGIC := '0';
	 SIGNAL MillisAlt : INTEGER;
	 SIGNAL SecondsAlt : INTEGER;
	 SIGNAL MinutesAlt : INTEGER;
	 SIGNAL startedAlt : STD_LOGIC := '0';
BEGIN

	 Timer_map: Timer PORT MAP(
        clock, started, Millis, Seconds, Minutes
    );
	 
	 TimerAlt_map: TimerAlt PORT MAP(
        clock, startedAlt, MillisAlt, SecondsAlt, MinutesAlt
    );
    
    servo_pwm1_map: servo_pwm1 PORT MAP(
        clock, reset, pos1, servo1
    );
	 
    servo_pwm2_map: servo_pwm2 PORT MAP(
        clock, reset, pos2, servo2
    );
	 
	 servo_pwm3_map: servo_pwm3 PORT MAP(
        clock, reset, pos3, servo3
    );
	 
	 servo_pwm4_map: servo_pwm4 PORT MAP(
        clock, reset, pos4, servo4
    );

    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,Ppad1_I,Button_1,Ppad2_I,Ppad3_I)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= State000;
            led9 <= '0';
            led8 <= '0';
            led7 <= '0';
            led6 <= '0';
            led5 <= '0';
            led4 <= '0';
            StateBit_1 <= '0';
            StateBit_2 <= '0';
            StateBit_3 <= '0';
			   pos2 <= 360;
	         pos1 <= 360;
				pos3 <= 360;
				pos4 <= 180;
				started <= '0';
				startedAlt <= '0';
				
        ELSE
            led9 <= '0';
            led8 <= '0';
            led7 <= '0';
            led6 <= '0';
            led5 <= '0';
            led4 <= '0';
            StateBit_1 <= '0';
            StateBit_2 <= '0';
            StateBit_3 <= '0';
				
            CASE fstate IS
                WHEN State000 =>
                    IF ((Ppad1_I = '1')) THEN
                        reg_fstate <= State001;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= State000;
                    END IF;
						  
						  started <= '0';
						  
						  startedAlt <= '0';

                    StateBit_3 <= '0';

                    led9 <= '1';

                    StateBit_2 <= '0';

                    StateBit_1 <= '0';
						  
						  pos1 <= 360;
						  pos2 <= 360;
						  pos3 <= 360;
						  pos4 <= 180; --start at final

						  
                WHEN State001 =>
                    IF ((Button_1 = '0')) THEN
                        reg_fstate <= State010;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= State001;
                    END IF;
						  
						  started <= '1';
						  
						  startedAlt <= '0';

                    StateBit_3 <= '1';

                    led8 <= '1';

                    StateBit_2 <= '0';

                    StateBit_1 <= '0';
						 
						  IF((Seconds >= 1 or Minutes > 0)) THEN
			           pos1 <= 50;
						  ELSE
						  pos1 <= 360;
						  pos3 <= 360;
						  END IF;

                WHEN State010 =>
                    IF ((Ppad2_I = '1')) THEN
                        reg_fstate <= State011;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= State010;
                    END IF;
						  
						  started <= '0';
						  
						  startedAlt <= '1';

                    StateBit_3 <= '0';

                    StateBit_2 <= '1';

                    StateBit_1 <= '0';

                    led7 <= '1';
						  
						  IF((SecondsAlt >= 2 or MinutesAlt > 0)) THEN
			           pos2 <= 0;
						  ELSE
						  pos2 <= 360;
						  pos3 <= 360;
						  END IF;
						  
                WHEN State011 =>
                    IF ((Ppad3_I = '1')) THEN
                        reg_fstate <= State100;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= State011;
                    END IF;
						  
						  startedAlt <= '0';
						  
						  started <= '1';

                    StateBit_3 <= '1';

                    StateBit_2 <= '1';

                    led6 <= '1';

                    StateBit_1 <= '0';
						  
						  IF((Seconds >= 1 or Minutes > 0)) THEN
			           pos3 <= 180;
						  pos4 <= 360;
						  ELSE
						  pos3 <= 360;
						  END IF;
						  
                WHEN State100 =>
                    IF ((Ppad2_I = '1')) THEN
                        reg_fstate <= State101;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= State100;
                    END IF;
						  
						  started <= '0';
						  
						  startedAlt <= '1';

                    led5 <= '1';

                    StateBit_3 <= '0';

                    StateBit_2 <= '0';

                    StateBit_1 <= '1';
						  
						  pos4 <= 360;
						  pos3 <= 180;
						  
						  
                WHEN State101 =>
                    IF ((Ppad3_I = '1')) THEN
                        reg_fstate <= State000;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= State101;
                    END IF;
						  
						  started <= '1';
						  
						  startedAlt <= '0';

                    led4 <= '1';

                    StateBit_3 <= '1';

                    StateBit_2 <= '0';

                    StateBit_1 <= '1';
						  
						  IF((Seconds >= 1 or Minutes > 0)) THEN
			           pos3 <= 0;
						  pos4 <= 180;	--**********
						  ELSE
						  pos3 <= 180;
						  END IF;
						  
                WHEN OTHERS => 
                    led9 <= 'X';
                    led8 <= 'X';
                    led7 <= 'X';
                    led6 <= 'X';
                    led5 <= 'X';
                    led4 <= 'X';
                    StateBit_1 <= 'X';
                    StateBit_2 <= 'X';
                    StateBit_3 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
